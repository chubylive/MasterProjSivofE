
`include "processing_element_if.sv"

package processing_element_test_pkg;

        `include "uvm_macros.svh"

        import uvm_pkg::*;

        `include "test_0.svh"

endpackage

